

module top (a, b, c, y);
input a, b, c;
output y;


xor (y, a, b, c);

endmodule
