
module top (a, b, c, y);
input a, b, c;
output y;


or (y, a, b, c);

endmodule
