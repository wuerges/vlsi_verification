module top (a, b, c, y);
input a, b, c;
output y;


and (y, a, b, c);

endmodule
